`timescale 1ns / 100ps

module tb_accumu_counter ();
	
	localparam CLK_PERIOD = 5;
	localparam SIZE = 3, NAME = "SCALE";
	localparam MAX_SIZE = SIZE - 1;
	localparam DEFAULT_SIZE = 3;

//Declare DUT signals
	integer tb_test_num;
	reg tb_clk;
	reg tb_n_rst;
	reg tb_clear;
	reg tb_count_enable;
	wire [MAX_SIZE:0] tb_count_out;
	wire tb_rollover_flag;

	//Declare under DUT
	reg [MAX_SIZE:0] expect_output;
	reg [MAX_SIZE:0] tb_test_data;
	reg expect_flag;

	always
	begin
		tb_clk = 1'b0;
		#(CLK_PERIOD/2.0);
		tb_clk = 1'b1;
		#(CLK_PERIOD/2.0);
	end


	accumu_counter DUT(.clk(tb_clk), .n_rst(tb_n_rst), .clear(tb_clear), .count_enable(tb_count_enable),.count_out(tb_count_out), .rollover_flag(tb_rollover_flag));

	initial
	begin
		//Initial all inputs
		tb_n_rst = 1'b0;
		tb_clear = 1'b0;
		tb_count_enable = 1'b1;
		tb_test_num = 0;
		tb_test_data = '0;
		expect_output = '0;
		expect_flag = 1'b0;

		#(0.1);

		//Test 1 check for proper reset
		@(negedge tb_clk);
		tb_test_num = tb_test_num + 1;
		tb_clear = 1'b0;
		tb_count_enable = 1'b0;
		@(posedge tb_clk);
		tb_n_rst = 1'b0;
		tb_test_data = '1;
		expect_output = '0;
		expect_flag = 0; 
		//@(posedge tb_clk);
		#1ns

		if ((expect_output == tb_count_out) && (expect_flag == tb_rollover_flag))
			$info("%s Case %0d:: PASSED", NAME, tb_test_num);
		else // Test case failed
			$error("%s Case %0d:: FAILED", NAME, tb_test_num);
		// De-assert reset for a cycle
		tb_n_rst = 1'b1;


		//Test 2 check for proper reset
		@(negedge tb_clk);
		tb_test_num = tb_test_num + 1;
		tb_clear = 1'b0;
		tb_count_enable = 1'b1;
		@(posedge tb_clk);	
		tb_n_rst = 1'b0;	
		tb_test_data = '1;
		expect_output = '0;
		expect_flag = 0;
		#1ns

		if ((expect_output == tb_count_out) && (expect_flag == tb_rollover_flag))
			$info("%s Case %0d:: PASSED", NAME, tb_test_num);
		else // Test case failed
			$error("%s Case %0d:: FAILED", NAME, tb_test_num);
		// De-assert reset for a cycle
		tb_n_rst <= 1'b1;


		//Test 3 check count enable
		@(negedge tb_clk);
		tb_test_num = tb_test_num + 1;
		tb_clear = 1'b0;
		tb_count_enable = 1'b1;
		@(posedge tb_clk);	
		tb_test_data = '0;
		expect_output = '0 + 1;
		expect_flag = 0;
		//@(posedge tb_clk);
		#1ns
		if ((expect_output == tb_count_out) && (expect_flag == tb_rollover_flag))
			$info("%s Case %0d:: PASSED", NAME, tb_test_num);
		else // Test case failed
			$error("%s Case %0d:: FAILED", NAME, tb_test_num);
		// De-assert reset for a cycle


		//Test 4 check count enable
		@(negedge tb_clk);
		tb_test_num = tb_test_num + 1;
		tb_clear = 1'b0;
		tb_count_enable = 1'b1;
		@(posedge tb_clk);	
		expect_output = 2;
		expect_flag = 1;
		//@(posedge tb_clk);
		#(1ns)
		
		if ((expect_output == tb_count_out) && (expect_flag == tb_rollover_flag))
			$info("%s Case %0d:: PASSED", NAME, tb_test_num);
		else // Test case failed
			$error("%s Case %0d:: FAILED", NAME, tb_test_num);
		// De-assert reset for a cycle
end
endmodule